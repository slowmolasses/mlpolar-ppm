// =============================================================================
// pkg_mlpolar.sv
// Package: Parameters for Multi-Level Polar Code over 1024-PPM Channel
//
// Channel model: 1024-ary PPM with transition matrix
//   P(l|k) = p         if l == k        (correct detection)
//          = q         if l == L+1      (erasure / photon lost)
//          = (1-p-q)/(L-1)  otherwise   (wrong slot / dark count)
//
// This implements the MLC-polar framework from Seidl et al. (2013):
//   - K=10 level sequential binary partition (SBP) lambda of the 1024-ary channel
//   - Each level i gets a polar component code of length N=256
//   - Component code rate R_i = I(B^i_lambda) (capacity rule, Sec. IV-A)
//   - Frozen set selected via BEC approximation to density evolution
//   - Multi-stage decoding (MSD): decoded level i feeds level i+1 as side info
//   - SP (natural binary) labeling: maximizes variance V_lambda(W) per Sec. IV-D
//
// Parameters tuned for: p=0.7, q=0.05, L=1024
// =============================================================================

package pkg_mlpolar;

  // -----------------------------------------------------------------------
  // Top-level dimensions
  // -----------------------------------------------------------------------
  localparam int L        = 1024;   // PPM alphabet size (# pulse slots)
  localparam int K_LEVELS = 10;     // log2(L) = number of SBP bit levels
  localparam int N        = 256;    // Component polar code block length
  localparam int LOG2N    = 8;      // n = log2(N), butterfly stages
  localparam int TOTAL_N  = K_LEVELS * N;  // 2560 total coded bits per block

  // -----------------------------------------------------------------------
  // Channel parameters (fixed-point approximations for FPGA arithmetic)
  // -----------------------------------------------------------------------
  // Represented as Q0.16 unsigned fixed-point (0..65535 = 0..1)
  localparam int FRAC_BITS = 16;
  localparam logic [FRAC_BITS-1:0] PROB_P = 16'hB333; // p=0.7
  localparam logic [FRAC_BITS-1:0] PROB_Q = 16'h0CCD; // q=0.05
  // r = (1-p-q)/(L-1) ≈ 2.444e-4 → 16-bit: ~16 (too small for Q0.16)
  // Use Q4.12 for r: 0.000244 * 4096 ≈ 1 → store as integer numerator
  // LLR computation handled in ppm_llr_compute with dedicated arithmetic

  // -----------------------------------------------------------------------
  // LLR quantization for SC decoder
  // -----------------------------------------------------------------------
  // LLRs are signed 8-bit: range [-128, 127], resolution 0.5 dB
  // Saturation at ±64 (6-bit useful range + saturation)
  localparam int LLR_BITS   = 8;
  localparam int LLR_MAX    =  64;
  localparam int LLR_MIN    = -64;
  typedef logic signed [LLR_BITS-1:0] llr_t;

  // -----------------------------------------------------------------------
  // Bit-level capacities I(B^i_lambda) for SP labeling, p=0.7, q=0.05
  // (computed offline by MLC bit-level mutual information decomposition)
  // Used to document frozen set selection; actual selection encoded in masks.
  // -----------------------------------------------------------------------
  // Level  0: I = 0.4160  ->  106 info bits, 150 frozen
  // Level  1: I = 0.5054  ->  129 info bits, 127 frozen
  // Level  2: I = 0.5740  ->  147 info bits, 109 frozen
  // Level  3: I = 0.6220  ->  159 info bits,  97 frozen
  // Level  4: I = 0.6532  ->  167 info bits,  89 frozen
  // Level  5: I = 0.6726  ->  172 info bits,  84 frozen
  // Level  6: I = 0.6842  ->  175 info bits,  81 frozen
  // Level  7: I = 0.6910  ->  177 info bits,  79 frozen
  // Level  8: I = 0.6949  ->  178 info bits,  78 frozen
  // Level  9: I = 0.6971  ->  178 info bits,  78 frozen
  // Total: 1588 info bits per block of 256 PPM symbols

  localparam int K_INFO [0:K_LEVELS-1] = '{106,129,147,159,167,172,175,177,178,178};

  // -----------------------------------------------------------------------
  // Frozen bit masks: FROZEN_MASK[level][i] = 1 iff channel i is frozen
  // 256-bit masks, one per bit level. Derived from BEC approximation.
  // Bit index i corresponds to synthetic polar channel B^(i)_{pi^n}.
  // Least significant bit = channel 0 (most unreliable → always frozen).
  // -----------------------------------------------------------------------
  // Each 256-bit value stored as four 64-bit hex words [255:192],[191:128],[127:64],[63:0]
  // NOTE: These masks are generated by scripts/mlpolar_design.py using exact
  // Bhattacharyya parameter density evolution (not the BEC approximation).
  // To regenerate: python scripts/mlpolar_design.py  and copy the printed block.
  localparam logic [255:0] FROZEN_MASK [0:K_LEVELS-1] = '{
    256'h000000000001011f0001037f177f7fff0017177f1fffffff7fffffffffffffff, // lvl 0
    256'h000000000000001700000117013f7fff0001037f177f7fff17ffffffffffffff, // lvl 1
    256'h00000000000000010000000701171fff00010117017f7fff177f7fffffffffff, // lvl 2
    256'h0000000000000001000000010017177f00000017011f7fff037f7fff7fffffff, // lvl 3
    256'h0000000000000001000000010003177f0000000701171fff013f7fff7fffffff, // lvl 4
    256'h0000000000000000000000010003077f00000007001717ff011f7fff7fffffff, // lvl 5
    256'h0000000000000000000000010001077f00000003001717ff011f3fff7fffffff, // lvl 6
    256'h0000000000000000000000010001037f00000003001717ff01173fff7fffffff, // lvl 7
    256'h0000000000000000000000010001037f00000003000717ff01173fff7fffffff, // lvl 8
    256'h0000000000000000000000010001037f00000003000717ff01173fff7fffffff  // lvl 9
  };

endpackage
